`default_nettype none

module myBigFSM
  (output logic [3:0] cMove,
   output logic win,
   output logic [15:0] hMove_all, cMove_all,
   input logic [3:0] hMove,
   input logic enter, clock, reset);

endmodule: myBigFSM